`timescale 1ns/1ps

module tb;

    // Testbench signals
    reg  [3:0] SW;
    reg        KEY;

    integer i;

    // DUT instantiation (edit name/ports if needed)
    // -----------------------------------------------
    // example:
    // my_module dut (
    //     .SW(SW),
    //     .KEY(KEY),
    //     .OUT(OUT)
    // );
    // -----------------------------------------------

    initial begin
        // Initialize
        SW  = 4'b0000;
        KEY = 1'b0;
        #5;

        // Test KEY = 0
        KEY = 1'b0;
        for (i = 0; i < 16; i = i + 1) begin
            SW = i[3:0];
            #5;
        end

        // Test KEY = 1
        KEY = 1'b1;
        for (i = 0; i < 16; i = i + 1) begin
            SW = i[3:0];
            #5;
        end

        // End simulation
        #10;
        $stop;
    end

endmodule
