// File Name: Selector.v
// Implements a 2-to-1 7-bit MUX
module Selector(
	input sel,            // Selector control input
	input [6:0] A, B,  // Selector data inputs
	output [6:0] F		  // Selector data outputs
	);
	

endmodule // Selector