// File Name: TestBench1.v
`timescale 1ns / 1ns
module TestBench1();
	reg [3:3] KEY;	// KEY = 0 --> SW[6:0],KEY = 1 --> SW[16:10]
	reg [17:0] SW;
	wire [6:0] LEDR;
	wire [6:0] HEX0;
	

	end
endmodule // TestBench1